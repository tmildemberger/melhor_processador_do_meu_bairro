library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity rom2 is
	port( 	clock				: in std_logic;
			endereco			: in unsigned(6 downto 0);
			dado				: out unsigned(17 downto 0)
	);
end entity;

architecture a_rom2 of rom2 is
	type mem is array(0 to 127) of unsigned(17 downto 0);
	constant conteudo_rom : mem := (
		0  => "011111101010101111",	-- MOV R7, #0x3f5   (0x3f5 tem o sinal extendido e se torna 0xfff5)
		1  => "110011010101111001",	-- MOV R6, #0x3579
		2  => "111111000011110000",	-- MOV R7, #0xf0f0
		3  => "011111101010101101",	-- MOV R5, #0x3f5   (0x3f5 tem o sinal extendido e se torna 0xfff5)
		4  => "001001101010111010",	-- MOV R2, #0x137
		5  => "000000101010000001",	-- MOV R1, #0x10
		6  => "000010101001101100", -- MOV R4, #77
		7  => "000000101000000011", -- MOV R3, #0
		8  => "101100010000110011", -- XOR R3, R6
		9  => "000000010100101110", -- SHL R6, #5
		10 => "101100000100001100", -- SUB R4, R1
		11 => "101100000000101101", -- ADD R5, R5
		12 => "101100000000001010", -- ADD R2, R1
		13 => "010001001100010111", -- OR  R7, #0x222   (0x222 tem o sinal extendido e se torna 0xfe22)
		14 => "000000011000011001", --ASHR R1, #3
		15 => "101100011100001111", -- ROL R7, R1
		16 => "001001100100011111", -- CMP R7, #0x123
		17 => "101100100100001100", -- CMP R4, R1
		18 => "101100101000111110", -- MOV R6, R7
		19 => "101100101000110101", -- MOV R5, R6
		20 => "000111101011011100",	-- MOV R4, #0xfb
		21 => "000000010101000100",	-- SHL R4, #8
		22 => "000110001101011100",	-- OR  R4, #0xcb
		23 => "101100101000000001",	-- MOV R1, R0
		24 => "000000000000000000", -- ADD R0, #0 (NOP)
		25 => "000000000000100001", -- ADD R1, #4
		26 => "101000000101100000", --JMPR UC, #5
		27 => "000000000000000000", -- 
		28 => "000000000000000000", -- 
		29 => "101011111111100000", --JMPR UC, #0xff
		30 => "000000000000000000", -- 
		31 => "101000011101000000", --JMPA UC, #0x1d
		32 => "101011111110100000", --JMPR UC, #0xfe
		33 => "000000000000000000", -- 
		34 => "000000000000000000",	-- 
		35 => "000000000000000000",	-- 
		36 => "000000000000000000", -- 
		37 => "000000000000000000", -- 
		38 => "000000000000000000", -- 
		39 => "000000000000000000", -- 
		40 => "000000000000000000", -- 
		41 => "000000000000000000", -- 
		42 => "000000000000000000", -- 
		43 => "000000000000000000", -- 
		44 => "000000000000000000", -- 
		45 => "000000000000000000", -- 
		46 => "000000000000000000",	-- 
		47 => "000000000000000000",	-- 
		48 => "000000000000000000",
		49 => "000000000000000000",
		others => (others => '0')
	);
	signal dado_interno			: unsigned(17 downto 0) := conteudo_rom(0);
begin
	process(clock)
	begin
		if (rising_edge(clock)) then
			dado_interno <= conteudo_rom(to_integer(endereco));
		end if;
	end process;
	
	dado <= dado_interno;
end architecture;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity rom_heap_sort is
	port( 	clock				: in std_logic;
			endereco			: in unsigned(6 downto 0);
			dado				: out unsigned(17 downto 0)
	);
end entity;

architecture a_rom_heap_sort of rom_heap_sort is
	type mem is array(0 to 127) of unsigned(17 downto 0);
	constant conteudo_rom : mem := (-- END. - INSTRUCAO
		0  => "101001001001010000",	-- 0x00 - CALLA UC, 0x49 - CALLA UC, fill_ram
		1  => "000000000000000000",	-- 0x01 - NOP
		2  => "101000001101010000",	-- 0x02 - CALLA UC, 0x0D - CALLA UC, heap_sort
		3  => "101011111111100000",	-- 0x03 - JMPR UC, 0xFF - JMPR UC, fim
		4  => "000000000100001100",	-- 0x04 - SUB  R4, #0x001
		5  => "000000011000001100",	-- 0x05 - ASHR R4, #0x001
		6  => "101111000000000000", -- 0x06 - RET
		7  => "000000010100001100", -- 0x07 - SHL  R4, #0x001
		8  => "000000000000001100", -- 0x08 - ADD  R4, #0x001
		9  => "101111000000000000", -- 0x09 - RET
		10 => "000000010100010100", -- 0x0A - SHL  R4, #0x001
		11 => "000000000000010100", -- 0x0B - ADD  R4, #0x002
		12 => "101111000000000000", -- 0x0C - RET
		13 => "101000010001110000", -- 0x0D - CALLR UC, 0x11 - CALLR UC, build_max_heap
		14 => "000000100100001111", -- 0x0E - CMP  R7, #0x001
		15 => "101000001110101111", -- 0x0F - JMPR ULE, 0x0E - JMPR UC, fim_heap_sort
		16 => "101100101000110101", -- 0x10 - MOV  R5, R6
		17 => "101100000000111101", -- 0x11 - ADD  R5, R7
		18 => "100011111111101011", -- 0x12 - MOV  R3, [R5 + #FF]
		19 => "100000000000110010", -- 0x13 - MOV  R2, [R6]
		20 => "100111111111101010",	-- 0x14 - MOV  [R5 + #FF], R2
		21 => "100100000000110011",	-- 0x15 - MOV  [R6], R3
		22 => "000000000100001111", -- 0x16 - SUB  R7, #0x001
		23 => "101100101000000100", -- 0x17 - MOV  R4, R0
		24 => "101110001100000101", -- 0x18 - PUSH R5
		25 => "101000101010010000", -- 0x19 - CALLA UC, 0x2A - CALLA UC, max_heapify
		26 => "101110000010000101", -- 0x1A - POP  R5
		27 => "000000000100001101", -- 0x1B - SUB  R5, #0x001
		28 => "000000100100001111", -- 0x1C - CMP  R7, #0x001
		29 => "101000010010001110", -- 0x1D - JMPA UGT, 0x12 - JMPA UGT, proximo_heap_sort
		30 => "101111000000000000", -- 0x1E - RET
		31 => "000000100100001111", -- 0x1F - CMP  R7, #0x001
		32 => "101000101001001111", -- 0x20 - JMPA ULE, 0x29 - JMPA ULE, fim_build_max_heap
		33 => "101100101000111100", -- 0x21 - MOV  R4, R7
		34 => "000000000100001100", -- 0x22 - SUB  R4, #0x001
		35 => "101011100000110000", -- 0x23 - CALLR UC, 0xE0 - CALLR UC, pai
		36 => "101110001100000100", -- 0x24 - PUSH R4
		37 => "101000101010010000", -- 0x25 - CALLA UC, 0x2A - CALLA UC, max_heapify
		38 => "101110000010000100", -- 0x26 - POP  R4
		39 => "000000000100001100", -- 0x27 - SUB  R4, #0x001
		40 => "101000100100000111", -- 0x28 - JMPA NN, 0x24 - JMPA NN, proximo_build_max_heap
		41 => "101111000000000000", -- 0x29 - RET
		42 => "101110001100000111", -- 0x2A - PUSH R7
		43 => "101110001100000110", -- 0x2B - PUSH R6
		44 => "000000000100001111", -- 0x2C - SUB  R7, #0x001
		45 => "101100101000110101", -- 0x2D - MOV  R5, R6
		46 => "101100000000100101", -- 0x2E - ADD  R5, R4
		47 => "100000000000101011", -- 0x2F - MOV  R3, [R5]
		48 => "101000000111010000", -- 0x30 - CALLA UC, 0x07 - CALLA UC, esquerda
		49 => "101100000000100110", -- 0x31 - ADD  R6, R4
		50 => "101100100100111100", -- 0x32 - CMP  R4, R7
		51 => "101000010001101110", -- 0x33 - JMPR UGT, 0x11 - JMPR UGT, nao_troca
		52 => "100000000000110010", -- 0x34 - MOV  R2, [R6]
		53 => "101000111100000010", -- 0x35 - JMPA EQ, 0x3C - JMPA EQ, pula_direita
		54 => "100000000001110001", -- 0x36 - MOV  R1, [R6 + #1]
		55 => "101100100100010001", -- 0x37 - CMP  R1, R2
		56 => "101000000011101111", -- 0x38 - JMPR ULE, 0x03 - JMPR ULE, pula_direita
		57 => "101100101000001010", -- 0x39 - MOV  R2, R1
		58 => "000000000000001110", -- 0x3A - ADD  R6, #1
		59 => "000000000000001100", -- 0x3B - ADD  R4, #1
		60 => "101100100100011010", -- 0x3C - CMP  R2, R3
		61 => "101001000101001111", -- 0x3D - JMPA ULE, 0x45 - JMPA ULE, nao_troca
		62 => "100100000000101010", -- 0x3E - MOV  [R5], R2
		63 => "101100101000110101", -- 0x3F - MOV  R5, R6
		64 => "101011000110110000", -- 0x40 - CALLR UC, 0xC6 - CALLR UC, esquerda
		65 => "101110000010000110", -- 0x41 - POP  R6
		66 => "101110001100000110", -- 0x42 - PUSH R6
		67 => "101100000000100110", -- 0x43 - ADD  R6, R4
		68 => "101000110010000000", -- 0x44 - JMPA UC, 0x32 - JMPA UC, volta
		69 => "100100000000101011", -- 0x45 - MOV  [R5], R3
		70 => "101110000010000110", -- 0x46 - POP  R6
		71 => "101110000010000111", -- 0x47 - POP  R7
		72 => "101111000000000000", -- 0x48 - RET
		73 => "110000000000100010", -- 0x49 - MOV  R6, #0x022
		74 => "000001101010010111", -- 0x4A - MOV  R7, #0x032
		75 => "000111101010000001", -- 0x4B - MOV  R1, #0x0F0
		76 => "000000010101000001", -- 0x4C - SHL  R1, #0x008
		77 => "000111001110000001", -- 0x4D - OR   R1, #0x0F0
		78 => "101100101000001010", -- 0x4E - MOV  R2, R1
		79 => "000000011000001001", -- 0x4F - ASHR R1, #0x001
		80 => "101100010000001010", -- 0x50 - XOR  R2, R1
		81 => "101100101000001011", -- 0x51 - MOV  R3, R1
		82 => "000000011000010011", -- 0x52 - ASHR R3, #0x002
		83 => "101100010000011010", -- 0x53 - XOR  R2, R3
		84 => "000000011001001011", -- 0x54 - ASHR R3, #0x009
		85 => "101100010000011010", -- 0x55 - XOR  R2, R3
		86 => "000000010000001010", -- 0x56 - XOR  R2, #0x001
		87 => "000000010101111010", -- 0x57 - SHL  R2, #0x00F
		88 => "101100010000010001", -- 0x58 - XOR  R1, R2
		89 => "101100101000001100", -- 0x59 - MOV  R4, R1
		90 => "101100101000001011", -- 0x5A - MOV  R3, R1
		91 => "000001001010000011", -- 0x5B - AND  R3, #0x020
		92 => "101000000001100010", -- 0x5C - JMPR Z, +1
		93 => "001011001011011100", -- 0x5D - AND  R4, #0x17B
		94 => "100100000000110100", -- 0x5E - MOV  [R6 + #0x00], R4
		95 => "000000000000001110", -- 0x5F - ADD  R6, #0x001
		96 => "000000000100001111", -- 0x60 - SUB  R7, #0x001
		97 => "101011101101100011", -- 0x61 - JMPR NZ, -19=0xED - JMPR NZ, voltafill_ram
		98 => "000001101000010110", -- 0x62 - MOV  R6, #0x022
		99 => "000001101010010111", -- 0x63 - MOV  R7, #0x032
		100 => "101111000000000000", -- 0x64 - RET
		others => (others => '0')
	);
	signal dado_interno			: unsigned(17 downto 0) := conteudo_rom(0);
begin
	process(clock)
	begin
		if (rising_edge(clock)) then
			dado_interno <= conteudo_rom(to_integer(endereco));
		end if;
	end process;
	
	dado <= dado_interno;
end architecture;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity rom_novos_formatos is
	port( 	clock				: in std_logic;
			endereco			: in unsigned(6 downto 0);
			dado				: out unsigned(17 downto 0)
	);
end entity;

architecture a_rom_novos_formatos of rom_novos_formatos is
	type mem is array(0 to 127) of unsigned(17 downto 0);
	constant conteudo_rom : mem := (-- END. - INSTRUÇÃO
		 0 => "000000000000000000", -- 0x00 - NOP
		 1 => "000000000000000000", -- 0x01 - NOP
		 2 => "000000000000000000", -- 0x02 - NOP
		 3 => "110000000000100010", -- 0x03 - MOV  R6, #0x022
		 4 => "000001101010010111", -- 0x04 - MOV  R7, #0x032
		 5 => "000111101010000001", -- 0x05 - MOV  R1, #0x0F0
		 6 => "000000010101000001", -- 0x06 - SHL  R1, #0x008
		 7 => "000111001110000001", -- 0x07 - OR   R1, #0x0F0
		 8 => "101100101000001010", -- 0x08 - MOV  R2, R1
		 9 => "000000011000001001", -- 0x09 - ASHR R1, #0x001
		10 => "101100010000001010", -- 0x0A - XOR  R2, R1
		11 => "101100101000001011", -- 0x0B - MOV  R3, R1
		12 => "000000011000010011", -- 0x0C - ASHR R3, #0x002
		13 => "101100010000011010", -- 0x0D - XOR  R2, R3
		14 => "000000011001001011", -- 0x0E - ASHR R3, #0x009
		15 => "101100010000011010", -- 0x0F - XOR  R2, R3
		16 => "000000010101111010", -- 0x10 - SHL  R2, #0x00F
		17 => "101100001100010001", -- 0x11 - OR   R1, R2
		18 => "101100101000001100", -- 0x12 - MOV  R4, R1
		19 => "101100101000001011", -- 0x13 - MOV  R3, R1
		20 => "000001001010000011", -- 0x14 - AND  R3, #0x020
		21 => "101000000001100010", -- 0x15 - JMPR Z, +1
		22 => "001011001011011100", -- 0x16 - AND  R4, #0x17B
		23 => "100100000000110100", -- 0x17 - MOV  [R6 + #0x00], R4
		24 => "000000000000001110", -- 0x18 - ADD  R6, #0x001
		25 => "000000000100001111", -- 0x19 - SUB  R7, #0x001
		26 => "101011101101100011", -- 0x1A - JMPR NZ, -19=0xED - JMPR NZ, volta_fill_ram
		27 => "000001101000010110", -- 0x1B - MOV  R6, #0x022
		28 => "000001101010010111", -- 0x1C - MOV  R7, #0x032
		29 => "000000000000000000", -- 0x1D - NOP
		30 => "110100011100101010", -- 0x1E - MOV  R6, #0x472A
		31 => "111111000011110000", -- 0x1F - MOV  R7, #0xF0F0
		32 => "101110001100000111", -- 0x20 - PUSH R7
		33 => "101110001100000110", -- 0x21 - PUSH R6
		34 => "101110000010000111", -- 0x22 - POP  R7
		35 => "101110000010000110", -- 0x23 - POP  R6
		36 => "101100101000111010", -- 0x24 - MOV  R2, R7
		37 => "101110001100000010", -- 0x25 - PUSH R2
		38 => "101110001100000100", -- 0x26 - PUSH R4
		39 => "101110100010000010", -- 0x27 - MOV  R2, SP
		40 => "000000000000001010", -- 0x28 - ADD  R2, #0x001
		41 => "101110100101000010", -- 0x29 - MOV  SP, R2
		42 => "101110000010000010", -- 0x2A - POP  R2
		43 => "101100100100111010", -- 0x2B - CMP  R2, R7
		44 => "101000101110010010", -- 0x2C - CALLA EQ, #0x2E
		45 => "101000000001100000", -- 0x2D - JMPR UC, #+1
		46 => "101111000000000000", -- 0x2E - RET
		47 => "100000010100110101", -- 0x2F - MOV  R5, [R6 + #0x14]
		48 => "101100010100110101", -- 0x30 - SHL  R5, R6
		49 => "101011111111100101", -- 0x31 - JMPR NV=0x5, #-1
		50 => "111100101011111110", -- 0x32 - MOV  R7, #0xCAFE
		51 => "000000101000101001", -- 0x33 - MOV  R1, #0x005
		52 => "101100100100001111", -- 0x34 - CMP  R7, R1
		53 => "101011111111101010", -- 0x35 - JMPR SGT=0xA, #-1
		54 => "101011111111101111", -- 0x36 - JMPR ULE=0xF, #-1
		55 => "101011111111100100", -- 0x37 - JMPR V=0x4, #-1
		56 => "101100101000111010", -- 0x38 - MOV  R2, R7
		57 => "101011111111101010", -- 0x39 - JMPR SGT=0xA, #-1
		58 => "101011111111101100", -- 0x3A - JMPR SLT=0xC, #-1
		59 => "101011111111101000", -- 0x3B - JMPR ULT=0x8, #-1
		60 => "101011111111101110", -- 0x3C - JMPR UGT=0xE, #-1
		61 => "101011111111100000", -- 0x3D - JMPR UC, #-1
		others => (others => '0')
	);
	signal dado_interno			: unsigned(17 downto 0) := conteudo_rom(0);
begin
	process(clock)
	begin
		if (rising_edge(clock)) then
			dado_interno <= conteudo_rom(to_integer(endereco));
		end if;
	end process;
	
	dado <= dado_interno;
end architecture;